class router_env extends uvm_env;

	// router reference
	router_reference reference;
	
	// router scoreboard
	router_scoreboard scoreboard;

	`uvm_component_utils_begin(router_env)
	`uvm_component_utils_end

	// UVM constructor
	function new(input string name, input uvm_component parent = null);
		super.new(name, parent);
	endfunction: new

	// UVM build_phase
	function void build_phase(uvm_phase phase);
		super.build_phase(phase);
		// instantiate the refrence model and scoreboard
		scoreboard = router_scoreboard::type_id::create("scoreboard", this);
		reference = router_reference::type_id::create("reference", this);
	endfunction: build_phase

	// UVM connect_phase
	function void connect_phase(uvm_phase phase);
		// connect the valid YAPP packet output port of the reference model to the input YAPP analysis imp of the scoreboard
		reference.sb_add_out.connect(scoreboard.sb_yapp_in);
	endfunction: connect_phase

endclass: router_env
